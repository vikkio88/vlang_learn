module console

import term

pub fn cls() {
	term.clear()
}
